`timescale 1ns / 1ps

module watch(
    input clk,
    input reset,
    input sec,
    input min,
    input hour,
    output [6:0] o_msec, 
    output [5:0] o_sec, o_min, 
    output [4:0] o_hour   
    );

    wire w_clk_100hz;                                                                                                                                                                                                                                                                                                                                                                                                                                         
    wire w_msec_tick, w_sec_tick, w_min_tick;

    clk_div_100hz_watch U_clk_div_100hz(
        .clk(clk),
        .reset(reset),
        .run(1'b1),                                       
        .o_clk(w_clk_100hz)
    );

    time_counter_watch #(.TICK_COUNT(100),.BIT_WIDTH(7)) U1_time_counter_msec(
        .clk(clk),
        .reset(reset),
        .tick(w_clk_100hz),
        .cnt(1'b0),
        .o_time(o_msec),
        .o_tick(w_msec_tick)
    );
                           
    time_counter_watch #(.TICK_COUNT(60),.BIT_WIDTH(6)) U2_time_counter_sec(
        .clk(clk),
        .reset(reset),
        .tick(w_msec_tick),
        .cnt(sec),
        .o_time(o_sec),
        .o_tick(w_sec_tick)
    );

    time_counter_watch #(.TICK_COUNT(60),.BIT_WIDTH(6)) U3_time_counter_min(
        .clk(clk),
        .reset(reset),
        .tick(w_sec_tick),
        .cnt(min),
        .o_time(o_min),
        .o_tick(w_min_tick)
    );

    time_counter_watch_hour #(.TICK_COUNT(24),.BIT_WIDTH(5)) U4_time_counter_hour(
        .clk(clk),
        .reset(reset),
        .tick(w_min_tick),
        .cnt(hour),
        .o_time(o_hour),
        .o_tick()
    );
endmodule

module clk_div_100hz_watch(
    input clk,
    input reset,
    input run,
    output o_clk
);

    parameter FCOUNT = 1_000_000; // 10 for debug
    reg [$clog2(FCOUNT) - 1 : 0] counter_reg, counter_next;
    reg clk_reg, clk_next;  
    assign o_clk = clk_reg;  // final output

    always @(posedge clk, posedge reset) begin
        if (reset) begin
            counter_reg <= 0;
            clk_reg <= 0;
        end
        else begin
            counter_reg <= counter_next;
            clk_reg <= clk_next;
        end
    end
// 
    always @(*) begin

        counter_next = counter_reg;
        clk_next = 1'b0;
        
        if(run == 1'b1) begin
            if (counter_reg == FCOUNT - 1) begin
                counter_next = 0;
                clk_next = 1'b1; 
            end 
            else begin
                counter_next = counter_reg + 1;
                clk_next = 1'b0;
            end
        end 
    end
endmodule

module time_counter_watch #(parameter TICK_COUNT = 100, BIT_WIDTH  = 7) (
    input clk,
    input reset,
    input tick,
    input cnt,  // cnt 입력 추가
    output [BIT_WIDTH - 1:0] o_time,
    output o_tick
);

    reg [$clog2(TICK_COUNT)-1:0] count_reg, count_next;
    reg tick_reg, tick_next;

    assign o_time = count_reg;
    assign o_tick = tick_reg;

    always @(posedge clk, posedge reset) begin
        if(reset) begin
            count_reg <= 0;
            tick_reg <=0;
        end 
        else begin
            count_reg <= count_next;
            tick_reg <= tick_next;
        end
    end

    // next logic
    always @(*) begin
        count_next = count_reg;
        tick_next = 1'b0; // tick_reg; 0 -> 1 -> 0
        
        // sec,min,hour 입력버튼 누르면 1 증가
        if(cnt == 1'b1) begin
            if (count_reg == TICK_COUNT - 1) begin
                count_next = 0;
                tick_next = 1'b1;
            end
            else begin
                count_next = count_reg + 1;
                tick_next = 1'b0;
            end
        end
        else if(tick == 1'b1) begin
            if (count_reg == TICK_COUNT - 1) begin
                count_next = 0;
                tick_next = 1'b1;
            end
            else begin
                count_next = count_reg + 1;
                tick_next = 1'b0;
            end
        end
    end
endmodule

module time_counter_watch_hour #(parameter TICK_COUNT = 24, BIT_WIDTH  = 5) (
    input clk,
    input reset,
    input tick,
    input cnt,  // cnt 입력 추가
    output [BIT_WIDTH - 1:0] o_time,
    output o_tick
);

    reg [$clog2(TICK_COUNT)-1:0] count_reg, count_next;
    reg tick_reg, tick_next;

    assign o_time = count_reg;
    assign o_tick = tick_reg;

    always @(posedge clk, posedge reset) begin
        if(reset) begin
            count_reg <= 12;
            tick_reg <=0;
        end 
        else begin
            count_reg <= count_next;
            tick_reg <= tick_next;
        end
    end

    // next logic
    always @(*) begin
        count_next = count_reg;
        tick_next = 1'b0; // tick_reg; 0 -> 1 -> 0
        
        // sec,min,hour 입력버튼 누르면 1 증가
        if(cnt == 1'b1) begin
            if (count_reg == TICK_COUNT - 1) begin
                count_next = 0;
                tick_next = 1'b1;
            end
            else begin
                count_next = count_reg + 1;
                tick_next = 1'b0;
            end
        end
        else if(tick == 1'b1) begin
            if (count_reg == TICK_COUNT - 1) begin
                count_next = 0;
                tick_next = 1'b1;
            end
            else begin
                count_next = count_reg + 1;
                tick_next = 1'b0;
            end
        end
    end
endmodule
`timescale 1ns / 1ns

module baud_tick_gen (
    input clk,
    input rst,
    output baud_tick
);

    parameter BAUD_RATE = 9600; //BAUD_RATE_19200 = 19200, ;
    localparam BAUD_COUNT = 100_000_000 / BAUD_RATE / 16;
    
    reg [$clog2(BAUD_COUNT)-1:0] cnt_reg, cnt_next;
    reg tick_reg, tick_next;

    assign baud_tick = tick_reg;

    always @(posedge clk, posedge rst) begin
        if(rst) begin
            tick_reg <= 0;
            cnt_reg <= 0;
        end
        else begin
            cnt_reg <= cnt_next;
            tick_reg <= tick_next;
        end 
    end

    always @(*) begin
        
       cnt_next = cnt_reg;
        tick_next = tick_reg;
        
        if(cnt_reg == BAUD_COUNT-1) begin
            cnt_next = 0;
            tick_next = 1'b1; 
        end
        else begin
            cnt_next = cnt_reg + 1;
            tick_next = 1'b0;
        end
    end
endmodule
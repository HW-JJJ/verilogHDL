`timescale 1ns / 1ps

module stopwatch_dp(
    input clk,
    input reset,
    input run,
    input clear,
    output [6:0] msec, sec, min, hour                
    );

    wire w_clk_100hz;
    wire w_msec_tick, w_sec_tick, w_min_tick;

    time_counter #(.TICK_COUNT(100)) U1_time_counter_msec(
        .clk(clk),
        .reset(reset),
        .tick(w_clk_100hz),
        .o_time(msec),
        .o_tick(w_msec_tick)
    );

    time_counter #(.TICK_COUNT(60)) U2_time_counter_sec(
        .clk(clk),
        .reset(reset),
        .tick(w_msec_tick),
        .o_time(sec),
        .o_tick(w_sec_tick)
    );

    time_counter #(.TICK_COUNT(60)) U3_time_counter_min(
        .clk(clk),
        .reset(reset),
        .tick(w_sec_tick),
        .o_time(min),
        .o_tick(w_min_tick)
    );

    time_counter #(.TICK_COUNT(24)) U4_time_counter_hour(
        .clk(clk),
        .reset(reset),
        .tick(w_min_tick),
        .o_time(hour),
        .o_tick()
    );

    clk_div_100hz U_clk_div_100hz(
        .clk(clk),
        .reset(reset),
        .run(run),
        .clear(clear),
        .o_clk(w_clk_100hz)
    );
endmodule

module clk_div_100hz(
    input clk,
    input reset,
    input run,
    input clear,
    output o_clk
);

    parameter FCOUNT = 10;
    reg [$clog2(FCOUNT) - 1 : 0] counter_reg, counter_next;
    reg clk_reg, clk_next;  // 출력을 f/f로 내보내기 위한
    
    assign o_clk = clk_reg;  // final output

    always @(posedge clk, posedge reset) begin
        if (reset) begin
            counter_reg <= 0;
            clk_reg <= 0;
        end
        else begin
            counter_reg <= counter_next;
            clk_reg <= clk_next;
        end
    end
// 
    always @(*) begin

        counter_next = counter_reg;
        clk_next = 1'b0;
        
        if(run == 1'b1) begin
            if (counter_reg == FCOUNT - 1) begin
                counter_next = 0;
                clk_next = 1'b1; // initial value
            end 
            else begin
                counter_next = counter_reg + 1;
                clk_next = 1'b0;
            end
        end 
        else if (clear == 1'b1) begin
            counter_next = 0;
            clk_next = 1'b0;
        end
    end
endmodule

module time_counter #(parameter TICK_COUNT = 100) (
    input clk,
    input reset,
    input tick,
    output [6:0] o_time,
    output o_tick
);

    reg [$clog2(TICK_COUNT)-1:0] count_reg, counter_next;
    reg tick_reg, tick_next;

    assign o_time = count_reg;
    assign o_tick = tick_reg;

    always @(posedge clk, posedge reset) begin
        if(reset) begin
            count_reg <= 0;
            tick_reg <=0;
        end 
        else begin
            count_reg <= counter_next;
            tick_reg <= tick_next;
        end
    end

    // next logic
    always @(*) begin

        counter_next = count_reg;
        tick_next = tick_reg;
        
        if(tick == 1'b1) begin
            if (count_reg == TICK_COUNT -1) begin
                counter_next = 0;
                tick_next = 1'b1;
            end
            else begin
                counter_next = count_reg + 1;
                tick_next = 1'b0;
            end
        end
    end


endmodule

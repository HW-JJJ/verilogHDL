`timescale 1ns / 1ps

module TOP_stopwatch(
    input clk,
    input reset,
    input btn_run,
    input btn_clear,
    output [6:0] o_msec, 
    output [5:0] o_sec, 
    output [5:0] o_min,
    output [4:0] o_hour
);
    wire w_run, w_clear;

    stopwatch_cu U_stopwatch_cu(
        .clk(clk),
        .reset(reset),
        .i_btn_run(btn_run),
        .i_btn_clear(btn_clear),
        .o_run(w_run),
        .o_clear(w_clear)
    );

    stopwatch_dp U_stopwatch_dp(
        .clk(clk),
        .reset(reset),
        .run(w_run),
        .clear(w_clear),
        .o_msec(o_msec),
        .o_sec(o_sec),
        .o_min(o_min),
        .o_hour(o_hour)                
    );
endmodule